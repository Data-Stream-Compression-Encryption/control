/*

Author: Alex Clarke
Date: 3/24/2015

This module tests the top level DSEC module

*/

module TB_DSEC;

reg clk;
reg rst;

reg key_config;
reg in_valid;
reg out_rcvd;
reg [63:0] data_in;

wire [63:0] data_out;
wire rdy, error, out_valid;

dsec u1(.clk(clk),.rst(rst),.data_in(data_in),.key_config(key_config),.in_valid(in_valid),.out_rcvd(out_rcvd),.rdy(rdy),.data_out(data_out),.error(error),.out_valid(out_valid));
 
// Generate a 50 MHz clock
initial
	clk = 1'b0;
always
	#10 clk = ~clk; 
	
initial begin
  rst = 1'b1;
  #20 rst = 1'b0;
  key_config = 1'b0;
  in_valid = 1'b0;
  out_rcvd = 1'b0;
  
  
  #20 key_config = 1'b1;
  data_in = 64'h9474B8E8C73BCA7D;
  #20 in_valid = 1'b1;
  #20 in_valid = 1'b0;
  data_in = 64'h8DA744E0C94E5E17;
  #20 in_valid = 1'b1;
  #20 in_valid = 1'b0;
  data_in = 64'h0CDB25E3BA3C6D79;
  #20 in_valid = 1'b1;
  #20 in_valid = 1'b0;
  key_config = 1'b0;
   
  data_in = 64'h9474B8E8C73BCA7D;
  #20 in_valid = 1'b1;
  #20 in_valid = 1'b0; 
  
  #20 out_rcvd = 1'b1;
  #20 out_rcvd = 1'b0;
  
  #20 key_config = 1'b1;
  data_in = 64'h0CDB25E3BA3C6D79;
  #20 in_valid = 1'b1;
  #20 in_valid = 1'b0;
  data_in = 64'h4784C4BA5006081F;
  #20 in_valid = 1'b1;
  #20 in_valid = 1'b0;
  data_in = 64'h1CF1FC126F2EF842;
  #20 in_valid = 1'b1;
  #20 in_valid = 1'b0;
  key_config = 1'b0;
   
  data_in = 64'h0CDB25E3BA3C6D79;
  #20 in_valid = 1'b1;
  #20 in_valid = 1'b0; 
	  
end



  
endmodule